library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity note2freq is
    port(
        midi_note : in unsigned(6 downto 0);
        rate : out signed(15 downto 0) -- basically frequency
    );
end note2freq;

architecture synth of note2freq is
    
begin
    with midi_note select rate <=
        16d"11" when 7d"0",
        16d"12" when 7d"1",
        16d"12" when 7d"2",
        16d"13" when 7d"3",
        16d"14" when 7d"4",
        16d"15" when 7d"5",
        16d"16" when 7d"6",
        16d"17" when 7d"7",
        16d"18" when 7d"8",
        16d"19" when 7d"9",
        16d"20" when 7d"10",
        16d"21" when 7d"11",
        16d"22" when 7d"12",
        16d"24" when 7d"13",
        16d"25" when 7d"14",
        16d"27" when 7d"15",
        16d"28" when 7d"16",
        16d"30" when 7d"17",
        16d"32" when 7d"18",
        16d"34" when 7d"19",
        16d"36" when 7d"20",
        16d"38" when 7d"21",
        16d"40" when 7d"22",
        16d"43" when 7d"23",
        16d"45" when 7d"24",
        16d"48" when 7d"25",
        16d"51" when 7d"26",
        16d"54" when 7d"27",
        16d"57" when 7d"28",
        16d"61" when 7d"29",
        16d"64" when 7d"30",
        16d"68" when 7d"31",
        16d"72" when 7d"32",
        16d"76" when 7d"33",
        16d"81" when 7d"34",
        16d"86" when 7d"35",
        16d"91" when 7d"36",
        16d"96" when 7d"37",
        16d"102" when 7d"38",
        16d"108" when 7d"39",
        16d"115" when 7d"40",
        16d"122" when 7d"41",
        16d"129" when 7d"42",
        16d"137" when 7d"43",
        16d"145" when 7d"44",
        16d"153" when 7d"45",
        16d"162" when 7d"46",
        16d"172" when 7d"47",
        16d"182" when 7d"48",
        16d"193" when 7d"49",
        16d"205" when 7d"50",
        16d"217" when 7d"51",
        16d"230" when 7d"52",
        16d"244" when 7d"53",
        16d"258" when 7d"54",
        16d"274" when 7d"55",
        16d"290" when 7d"56",
        16d"307" when 7d"57",
        16d"325" when 7d"58",
        16d"345" when 7d"59",
        16d"365" when 7d"60",
        16d"387" when 7d"61",
        16d"410" when 7d"62",
        16d"434" when 7d"63",
        16d"460" when 7d"64",
        16d"488" when 7d"65",
        16d"517" when 7d"66",
        16d"548" when 7d"67",
        16d"580" when 7d"68",
        16d"615" when 7d"69",
        16d"651" when 7d"70",
        16d"690" when 7d"71",
        16d"731" when 7d"72",
        16d"775" when 7d"73",
        16d"821" when 7d"74",
        16d"869" when 7d"75",
        16d"921" when 7d"76",
        16d"976" when 7d"77",
        16d"1034" when 7d"78",
        16d"1096" when 7d"79",
        16d"1161" when 7d"80",
        16d"1230" when 7d"81",
        16d"1303" when 7d"82",
        16d"1380" when 7d"83",
        16d"1463" when 7d"84",
        16d"1550" when 7d"85",
        16d"1642" when 7d"86",
        16d"1739" when 7d"87",
        16d"1843" when 7d"88",
        16d"1953" when 7d"89",
        16d"2069" when 7d"90",
        16d"2192" when 7d"91",
        16d"2322" when 7d"92",
        16d"2460" when 7d"93",
        16d"2606" when 7d"94",
        16d"2761" when 7d"95",
        16d"2926" when 7d"96",
        16d"3100" when 7d"97",
        16d"3284" when 7d"98",
        16d"3479" when 7d"99",
        16d"3686" when 7d"100",
        16d"3906" when 7d"101",
        16d"4138" when 7d"102",
        16d"4384" when 7d"103",
        16d"4645" when 7d"104",
        16d"4921" when 7d"105",
        16d"5213" when 7d"106",
        16d"5523" when 7d"107",
        16d"5852" when 7d"108",
        16d"6200" when 7d"109",
        16d"6569" when 7d"110",
        16d"6959" when 7d"111",
        16d"7373" when 7d"112",
        16d"7812" when 7d"113",
        16d"8276" when 7d"114",
        16d"8768" when 7d"115",
        16d"9290" when 7d"116",
        16d"9842" when 7d"117",
        16d"10427" when 7d"118",
        16d"11047" when 7d"119",
        16d"11704" when 7d"120",
        16d"12400" when 7d"121",
        16d"13138" when 7d"122",
        16d"13919" when 7d"123",
        16d"14747" when 7d"124",
        16d"15624" when 7d"125",
        16d"16553" when 7d"126",
        16d"17537" when 7d"127",
        16d"0" when others;
end;
